/**
  *   NOTE THAT THIS IS DRIVING THE SPI SLAVE
  */

interface gr_spi_if(input clk, input reset);
  
  logic   ss;
  logic   sclk;
  logic   mosi;
  logic   miso;

  
endinterface
